`timescale 1ns / 1ps

module IIR_fold(
clk,
rst,
a,b,c,d,
x,
y
);

input clk,rst;
input[7:0] a,b,c,d;
input[7:0] x;
output[7:0] y;

/*************** Your code here ***************/



/********************* Done *********************/

endmodule
